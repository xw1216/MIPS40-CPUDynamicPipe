`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 
// Create Date: 2021/11/03 11:24:14
// Design Name: 
// Module Name: UEXT16
// 
//////////////////////////////////////////////////////////////////////////////////


module uext16
(
    input  wire [15:0] din,
    output wire [31:0] dout
);

assign dout = { 16'b0, din[15:0]}; 
endmodule
