`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 
// Create Date: 2021/11/04 12:02:02
// Design Name: 
// Module Name: EXT18
// 
//////////////////////////////////////////////////////////////////////////////////


module ext18
(
    input  wire [15:0] din,
    output wire [31:0] dout
);


assign dout = { {14{din[15]}}, din[15:0], 2'b00 };

endmodule
