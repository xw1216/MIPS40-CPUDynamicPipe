`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 
// Create Date: 2021/11/03 11:24:14
// Design Name: 
// Module Name: EXT16
// 
//////////////////////////////////////////////////////////////////////////////////


module ext16
(
    input  wire [15:0] din,
    output wire [31:0] dout
);

assign dout = { {16{din[15]}}, din[15:0]}; 
endmodule
